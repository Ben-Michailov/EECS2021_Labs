module labM;
wire [31:0] rd1, rd2;
reg clk, w, flag;
reg [31:0] wd;
reg[4:0] rs1, rs2, wn;
integer i;
rf myRF(rd1, rd2, rs1, rs2, wn, wd, clk, w);
initial
begin
    flag = $value$plusargs("w=%b", w);
    for (i = 0; i < 32; i = i + 1)
    begin
        clk = 0;
        wd = i * i;
        wn = i;
        clk = 1;
        #1;
    end

    repeat(10)
    begin
        rs1 = $random;
        rs2 = $random;
        #1
        $display("clk=%b, w=%b, rs1=%d, rs2=%d, rd1=%d, rd2=%d", clk,w, rs1, rs2, rd1, rd2);

    end

    $finish;
end

endmodule